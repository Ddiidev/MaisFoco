module contact

import veb
import mf_core.logger

pub struct ContactController {
	veb.Context
pub:
	log logger.ILogger
}
