module contact

import veb
import shareds.logger

pub struct ContactController {
	veb.Context
pub:
	log logger.ILogger
}
