module home

import veb
import mf_core.logger

pub struct HomePage {
	veb.Controller
pub mut:
	log logger.ILogger
}
