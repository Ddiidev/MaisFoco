module about

import veb
import mf_core.logger

pub struct AboutCrontoller {
	veb.Context
pub:
	log logger.ILogger
}
