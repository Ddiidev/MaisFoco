module about

import veb
import shareds.logger

pub struct AboutCrontoller {
	veb.Context
pub:
	log logger.ILogger
}
